
ENTITY top_level_blk_mem_gen_0_0 IS
  PORT (
    clka : IN STD_LOGIC;
    addra : IN STD_LOGIC_VECTOR(13 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END top_level_blk_mem_gen_0_0;
  
  
  
  
